library verilog;
use verilog.vl_types.all;
entity altera_tristate_controller_aggregator is
    generic(
        AV_ADDRESS_W    : integer := 32;
        AV_DATA_W       : integer := 32;
        AV_BYTEENABLE_W : integer := 4
    );
    port(
        av_address      : in     vl_logic_vector;
        av_read         : in     vl_logic;
        av_write        : in     vl_logic;
        av_byteenable   : in     vl_logic_vector;
        av_writebyteenable: in     vl_logic_vector;
        av_readdata     : out    vl_logic_vector;
        av_writedata    : in     vl_logic_vector;
        av_lock         : in     vl_logic;
        av_chipselect   : in     vl_logic;
        av_outputenable : in     vl_logic;
        av_waitrequest  : out    vl_logic;
        av_begintransfer: in     vl_logic;
        tcm0_request    : out    vl_logic;
        tcm0_grant      : in     vl_logic;
        tcm0_address    : out    vl_logic_vector;
        tcm0_read       : out    vl_logic;
        tcm0_read_n     : out    vl_logic;
        tcm0_write      : out    vl_logic;
        tcm0_write_n    : out    vl_logic;
        tcm0_begintransfer: out    vl_logic;
        tcm0_begintransfer_n: out    vl_logic;
        tcm0_byteenable : out    vl_logic_vector;
        tcm0_byteenable_n: out    vl_logic_vector;
        tcm0_writedata  : out    vl_logic_vector;
        tcm0_readdata   : in     vl_logic_vector;
        tcm0_data_outen : out    vl_logic;
        tcm0_writebyteenable: out    vl_logic_vector;
        tcm0_writebyteenable_n: out    vl_logic_vector;
        tcm0_outputenable: out    vl_logic;
        tcm0_outputenable_n: out    vl_logic;
        tcm0_chipselect : out    vl_logic;
        tcm0_chipselect_n: out    vl_logic;
        tcm0_waitrequest: in     vl_logic;
        tcm0_waitrequest_n: in     vl_logic;
        tcm0_lock       : out    vl_logic;
        tcm0_lock_n     : out    vl_logic;
        tcm0_resetrequest: in     vl_logic;
        tcm0_resetrequest_n: in     vl_logic;
        tcm0_irq_in     : in     vl_logic;
        tcm0_irq_in_n   : in     vl_logic;
        tcm0_reset_output: out    vl_logic;
        tcm0_reset_output_n: out    vl_logic;
        c0_request      : in     vl_logic;
        c0_grant        : out    vl_logic;
        c0_uav_write    : in     vl_logic;
        irq_out         : out    vl_logic;
        reset_out       : out    vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AV_ADDRESS_W : constant is 1;
    attribute mti_svvh_generic_type of AV_DATA_W : constant is 1;
    attribute mti_svvh_generic_type of AV_BYTEENABLE_W : constant is 1;
end altera_tristate_controller_aggregator;
