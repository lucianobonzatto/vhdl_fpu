library verilog;
use verilog.vl_types.all;
entity system_0 is
    port(
        clk_50          : in     vl_logic;
        bidir_port_to_and_from_the_SD_DAT: inout  vl_logic;
        out_port_from_the_led_red: out    vl_logic_vector(17 downto 0);
        zs_addr_from_the_sdram_0: out    vl_logic_vector(11 downto 0);
        zs_ba_from_the_sdram_0: out    vl_logic_vector(1 downto 0);
        zs_cas_n_from_the_sdram_0: out    vl_logic;
        zs_cke_from_the_sdram_0: out    vl_logic;
        zs_cs_n_from_the_sdram_0: out    vl_logic;
        zs_dq_to_and_from_the_sdram_0: inout  vl_logic_vector(15 downto 0);
        zs_dqm_from_the_sdram_0: out    vl_logic_vector(1 downto 0);
        zs_ras_n_from_the_sdram_0: out    vl_logic;
        zs_we_n_from_the_sdram_0: out    vl_logic;
        tri_state_bridge_0_data: inout  vl_logic_vector(7 downto 0);
        tri_state_bridge_0_readn: out    vl_logic_vector(0 downto 0);
        write_n_to_the_cfi_flash_0: out    vl_logic_vector(0 downto 0);
        tri_state_bridge_0_address: out    vl_logic_vector(21 downto 0);
        select_n_to_the_cfi_flash_0: out    vl_logic_vector(0 downto 0);
        reset_n         : in     vl_logic;
        bidir_port_to_and_from_the_SD_CMD: inout  vl_logic;
        in_port_to_the_button_pio: in     vl_logic_vector(3 downto 0);
        USB_DATA_to_and_from_the_ISP1362: inout  vl_logic_vector(15 downto 0);
        USB_ADDR_from_the_ISP1362: out    vl_logic_vector(1 downto 0);
        USB_RD_N_from_the_ISP1362: out    vl_logic;
        USB_WR_N_from_the_ISP1362: out    vl_logic;
        USB_CS_N_from_the_ISP1362: out    vl_logic;
        USB_RST_N_from_the_ISP1362: out    vl_logic;
        USB_INT0_to_the_ISP1362: in     vl_logic;
        USB_INT1_to_the_ISP1362: in     vl_logic;
        out_port_from_the_SD_CLK: out    vl_logic;
        out_port_from_the_led_green: out    vl_logic_vector(8 downto 0);
        in_port_to_the_switch_pio: in     vl_logic_vector(17 downto 0);
        LCD_RS_from_the_lcd_16207_0: out    vl_logic;
        LCD_RW_from_the_lcd_16207_0: out    vl_logic;
        LCD_data_to_and_from_the_lcd_16207_0: inout  vl_logic_vector(7 downto 0);
        LCD_E_from_the_lcd_16207_0: out    vl_logic;
        rxd_to_the_uart_0: in     vl_logic;
        txd_from_the_uart_0: out    vl_logic;
        audio_0_oAUD_DATA: out    vl_logic;
        audio_0_oAUD_LRCK: out    vl_logic;
        audio_0_oAUD_BCK: out    vl_logic;
        audio_0_oAUD_XCK: out    vl_logic;
        audio_0_iCLK_18_4: in     vl_logic;
        vga_0_VGA_R     : out    vl_logic_vector(9 downto 0);
        vga_0_VGA_G     : out    vl_logic_vector(9 downto 0);
        vga_0_VGA_B     : out    vl_logic_vector(9 downto 0);
        vga_0_VGA_HS    : out    vl_logic;
        vga_0_VGA_VS    : out    vl_logic;
        vga_0_VGA_SYNC  : out    vl_logic;
        vga_0_VGA_BLANK : out    vl_logic;
        vga_0_VGA_CLK   : out    vl_logic;
        vga_0_iCLK_25   : in     vl_logic;
        dm9000a_iOSC_50 : in     vl_logic;
        dm9000a_ENET_DATA: inout  vl_logic_vector(15 downto 0);
        dm9000a_ENET_CMD: out    vl_logic;
        dm9000a_ENET_RD_N: out    vl_logic;
        dm9000a_ENET_WR_N: out    vl_logic;
        dm9000a_ENET_CS_N: out    vl_logic;
        dm9000a_ENET_RST_N: out    vl_logic;
        dm9000a_ENET_CLK: out    vl_logic;
        dm9000a_ENET_INT: in     vl_logic;
        seg7_display_oSEG0: out    vl_logic_vector(6 downto 0);
        seg7_display_oSEG1: out    vl_logic_vector(6 downto 0);
        seg7_display_oSEG2: out    vl_logic_vector(6 downto 0);
        seg7_display_oSEG3: out    vl_logic_vector(6 downto 0);
        seg7_display_oSEG4: out    vl_logic_vector(6 downto 0);
        seg7_display_oSEG5: out    vl_logic_vector(6 downto 0);
        seg7_display_oSEG6: out    vl_logic_vector(6 downto 0);
        seg7_display_oSEG7: out    vl_logic_vector(6 downto 0);
        sram_0_avalon_slave_0_export_DQ: inout  vl_logic_vector(15 downto 0);
        sram_0_avalon_slave_0_export_ADDR: out    vl_logic_vector(17 downto 0);
        sram_0_avalon_slave_0_export_UB_N: out    vl_logic;
        sram_0_avalon_slave_0_export_LB_N: out    vl_logic;
        sram_0_avalon_slave_0_export_WE_N: out    vl_logic;
        sram_0_avalon_slave_0_export_CE_N: out    vl_logic;
        sram_0_avalon_slave_0_export_OE_N: out    vl_logic
    );
end system_0;
