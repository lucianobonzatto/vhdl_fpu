library verilog;
use verilog.vl_types.all;
entity tornado_system_0_epcs_controller_atom is
    port(
        dclkin          : in     vl_logic;
        oe              : in     vl_logic;
        scein           : in     vl_logic;
        sdoin           : in     vl_logic;
        data0out        : out    vl_logic
    );
end tornado_system_0_epcs_controller_atom;
